`define HASTI_TRANS_IDLE 2'b00
`define HASTI_TRANS_BUSY 2'b01
`define HASTI_TRANS_NONSEQ 2'b10
`define HASTI_TRANS_SEQ 2'b11

`define HASTI_BURST_SINGLE 3'b0

`define HASTI_MASTER_NO_LOCK 1'b0

`define HASTI_RESP_OKAY 1'b0
`define HASTI_RESP_ERROR 1'b1

