`define RV32_LOAD     0000011
`define RV32_STORE    0100011
`define RV32_MADD     1000011
`define RV32_BRANCH   1100011

`define RV32_LOAD_FP  0000111
`define RV32_STORE_FP 0100111 
`define RV32_MSUB     1000111
`define RV32_JALR     1100111

`define RV32_CUSTOM_0 0001011
`define RV32_CUSTOM_1 0101011
`define RV32_NMSUB    1001011
// 1101011 is reserved

`define RV32_MISC_MEM 0001111
`define RV32_AMO      0101111
`define RV32_NMADD    1001111
`define RV32_JAL      1101111

`define RV32_OP_IMM   0010011
`define RV32_OP       0110011
`define RV32_OP_FP    1010011
`define RV32_SYSTEM   1110011

`define RV32_AUIPC    0010111
`define RV32_LUI      0110111
// 1010111 is reserved
// 1110111 is reserved

// 0011011 is RV64-specific
// 0111011 is RV64-specific
`define RV32_CUSTOM_2 1011011
`define RV32_CUSTOM_3 1111011
