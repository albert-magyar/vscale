`define HASTI_TRANS_IDLE 2'b00
`define HASTI_TRANS_BUSY 2'b01
`define HASTI_TRANS_NONSEQ 2'b10
`define HASTI_TRANS_SEQ 2'b11

`define HASTI_NO_PROT 4'b0

`define HASTI_BURST_SINGLE 3'b0

`define HASTI_MASTER_NO_LOCK 1'b0

`define HASTI_RESP_OKAY 1'b0
`define HASTI_RESP_ERROR 1'b1

`define HASTI_SIZE_BYTE     3'b000
`define HASTI_SIZE_HALFWORD 3'b001
`define HASTI_SIZE_WORD     3'b010
