`define ALU_OP_ADD  0
`define ALU_OP_SL   1
`define ALU_OP_XOR  4
`define ALU_OP_OR   6
`define ALU_OP_AND  7
`define ALU_OP_SR   5
`define ALU_OP_SEQ  8
`define ALU_OP_SNE  9
`define ALU_OP_SUB  10
`define ALU_OP_SRA  11
`define ALU_OP_SLT  12
`define ALU_OP_SGE  13
`define ALU_OP_SLTU 14
`define ALU_OP_SGEU 15
